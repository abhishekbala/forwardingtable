library verilog;
use verilog.vl_types.all;
entity entity_table_vlg_vec_tst is
end entity_table_vlg_vec_tst;

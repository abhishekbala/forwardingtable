library verilog;
use verilog.vl_types.all;
entity camTestBench_vlg_vec_tst is
end camTestBench_vlg_vec_tst;

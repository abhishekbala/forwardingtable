library verilog;
use verilog.vl_types.all;
entity fwdTable_vlg_vec_tst is
end fwdTable_vlg_vec_tst;
